module cube532
(
  input clk,
  input  [7:0]  in,
  output [23:0] out
);

// Your Code Here

endmodule
