`timescale 1ns / 1ps

module mask532
(
  input [4:0] 	n,
  input [31:0]  value_in,
  output [31:0] value_out
);

	// Your Code Here

endmodule